library verilog;
use verilog.vl_types.all;
entity openmips_min_sopc is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic
    );
end openmips_min_sopc;
