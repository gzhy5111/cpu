library verilog;
use verilog.vl_types.all;
entity openmips_min_sopc_tb is
end openmips_min_sopc_tb;
